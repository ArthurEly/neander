library verilog;
use verilog.vl_types.all;
entity ulaoitobits_vlg_vec_tst is
end ulaoitobits_vlg_vec_tst;
