library verilog;
use verilog.vl_types.all;
entity decodneanderinstructions_vlg_vec_tst is
end decodneanderinstructions_vlg_vec_tst;
