library verilog;
use verilog.vl_types.all;
entity registradoroitobits_vlg_vec_tst is
end registradoroitobits_vlg_vec_tst;
