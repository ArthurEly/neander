library verilog;
use verilog.vl_types.all;
entity registradordoisbits_vlg_check_tst is
    port(
        N_out           : in     vl_logic;
        Z_out           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end registradordoisbits_vlg_check_tst;
