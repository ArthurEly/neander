library verilog;
use verilog.vl_types.all;
entity lab041_vlg_vec_tst is
end lab041_vlg_vec_tst;
