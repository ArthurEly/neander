library verilog;
use verilog.vl_types.all;
entity ulaumbit_vlg_vec_tst is
end ulaumbit_vlg_vec_tst;
