library verilog;
use verilog.vl_types.all;
entity ulaumbit_vlg_check_tst is
    port(
        cout            : in     vl_logic;
        \out\           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ulaumbit_vlg_check_tst;
