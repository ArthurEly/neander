library verilog;
use verilog.vl_types.all;
entity registradordoisbits_vlg_vec_tst is
end registradordoisbits_vlg_vec_tst;
