library verilog;
use verilog.vl_types.all;
entity acumuladorumbit_vlg_vec_tst is
end acumuladorumbit_vlg_vec_tst;
