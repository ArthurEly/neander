library verilog;
use verilog.vl_types.all;
entity parteoperativa_vlg_vec_tst is
end parteoperativa_vlg_vec_tst;
