library verilog;
use verilog.vl_types.all;
entity lab041 is
    port(
        d3              : out    vl_logic;
        v               : in     vl_logic;
        a1              : in     vl_logic;
        a0              : in     vl_logic;
        d2              : out    vl_logic;
        d1              : out    vl_logic;
        d0              : out    vl_logic
    );
end lab041;
