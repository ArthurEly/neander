library verilog;
use verilog.vl_types.all;
entity contadortresbits_vlg_check_tst is
    port(
        a0              : in     vl_logic;
        a1              : in     vl_logic;
        a2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end contadortresbits_vlg_check_tst;
