library verilog;
use verilog.vl_types.all;
entity partedecontrole_vlg_vec_tst is
end partedecontrole_vlg_vec_tst;
