library verilog;
use verilog.vl_types.all;
entity acumulador_vlg_vec_tst is
end acumulador_vlg_vec_tst;
