library verilog;
use verilog.vl_types.all;
entity \lab041-bkp\ is
    port(
        d15             : out    vl_logic;
        a3              : in     vl_logic;
        a2              : in     vl_logic;
        d14             : out    vl_logic;
        d13             : out    vl_logic;
        d12             : out    vl_logic;
        d11             : out    vl_logic;
        a1b             : in     vl_logic;
        a0b             : in     vl_logic;
        d10             : out    vl_logic;
        d9              : out    vl_logic;
        d8              : out    vl_logic
    );
end \lab041-bkp\;
