library verilog;
use verilog.vl_types.all;
entity lab0412_vlg_vec_tst is
end lab0412_vlg_vec_tst;
