library verilog;
use verilog.vl_types.all;
entity lab041_vlg_check_tst is
    port(
        d0              : in     vl_logic;
        d1              : in     vl_logic;
        d2              : in     vl_logic;
        d3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab041_vlg_check_tst;
