library verilog;
use verilog.vl_types.all;
entity pcumbit_vlg_vec_tst is
end pcumbit_vlg_vec_tst;
