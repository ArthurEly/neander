library verilog;
use verilog.vl_types.all;
entity contadortresbits_vlg_vec_tst is
end contadortresbits_vlg_vec_tst;
