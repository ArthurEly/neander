library verilog;
use verilog.vl_types.all;
entity uc_vlg_vec_tst is
end uc_vlg_vec_tst;
