library verilog;
use verilog.vl_types.all;
entity decodula_vlg_vec_tst is
end decodula_vlg_vec_tst;
