library verilog;
use verilog.vl_types.all;
entity lab0412_vlg_check_tst is
    port(
        d0              : in     vl_logic;
        d1              : in     vl_logic;
        d2              : in     vl_logic;
        d3              : in     vl_logic;
        d4              : in     vl_logic;
        d5              : in     vl_logic;
        d6              : in     vl_logic;
        d7              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab0412_vlg_check_tst;
