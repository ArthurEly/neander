library verilog;
use verilog.vl_types.all;
entity decod3x8 is
    port(
        d3              : out    vl_logic;
        a2              : in     vl_logic;
        a1              : in     vl_logic;
        a0              : in     vl_logic;
        d2              : out    vl_logic;
        d1              : out    vl_logic;
        d0              : out    vl_logic;
        d7              : out    vl_logic;
        d6              : out    vl_logic;
        d5              : out    vl_logic;
        d4              : out    vl_logic
    );
end decod3x8;
